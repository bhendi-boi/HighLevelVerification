
interface intf (
    input logic clk,
    reset
);

  //declaring the signals

  logic [3:0] a;
  logic [3:0] b;
  logic add_sub;
  logic [6:0] cout;

endinterface
