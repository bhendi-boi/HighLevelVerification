module ahb_slave (
    ahb_if ahb_bus
);
  // DUMMY SLAVE
endmodule

