module env (
    input reset,
    input txclk,
    input ld_tx_data,
    input [7:0] tx_data,
    input tx_enable,
    input tx_out,
    input tx_empty,
    input rxclk,
    input uld_rx_data,
    input [7:0] rx_data,
    input rx_enable,
    input rx_in,
    input rx_empty,
);

  

endmodule
