
//gets the packet from generator and drive the transaction paket items into interface (interface is connected to DUT, so the items driven into interface signal will get driven in to DUT) 

class driver;

  //used to count the number of transactions
  int no_transactions;

  //creating virtual interface handle
  virtual counter_inf vif;

  //creating mailbox handle
  mailbox gen2driv;

  //constructor
  function new(virtual counter_inf vif, mailbox gen2driv);
    //getting the interface
    this.vif = vif;
    //getting the mailbox handles from  environment 
    this.gen2driv = gen2driv;
  endfunction

  //Reset task, Reset the Interface signals to default/initial values
  task reset;
    wait (vif.rst);
    $display("[ DRIVER ] ----- Reset Started -----");
    vif.load <= 1;
    vif.data_in <= 0;
    wait (!vif.rst);
    $display("[ DRIVER ] ----- Reset Ended   -----");
  endtask

  //drivers the transaction items to interface signals
  task main;
    forever begin
      transaction trans;
      gen2driv.get(trans);
      //@(posedge vif.clk);

      vif.load    <= trans.load;
      vif.data_in <= trans.data_in;
      vif.up_down <= trans.up_down;
      @(posedge vif.clk);

      trans.data_out = vif.data_out;
      //@(posedge vif.clk);
      trans.display("[ Driver ]");
      no_transactions++;
    end
  endtask

endclass
