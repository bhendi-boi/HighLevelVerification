package automatic my_package;
    class MemTrans;
        bit [7:0] data_in;
        bit [3:0] address;
        Statistics stats;
        function new();
            data_in = 3;
            address Si
            stats = new();
        endfunction

        function copy();
                        
        endfunction
    endclass;
endpackage