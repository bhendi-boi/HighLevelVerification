
`include "environment.sv"

program test (
    counter_inf i_intf
);

  class my_trans extends transaction;

    function void pre_randomize();
      load.rand_mode(0);
      data_in.rand_mode(0);

      load = 1;
      data_in = 12;

    endfunction

  endclass

  //declaring environment instance
  environment env;
  my_trans my_tr;

  initial begin
    //creating environment
    env = new(i_intf);

    my_tr = new();

    //setting the repeat count of generator as 4, means to generate 4 packets
    env.gen.repeat_count = 4;

    env.gen.trans = my_tr;

    //calling run of env, it interns calls generator and driver main tasks.
    my_tr.pre_randomize();
    env.run();
  end
endprogram
